// $Id: $
// File name:   USB_tx_top_level.sv
// Created:     12/1/2017
// Author:      Michael Toner
// Lab Section: 337-05
// Version:     1.0  Initial Design Entry
// Description: Top level module for transmitting USB module .
