// $Id: $
// File name:   tb_helper.sv
// Created:     12/6/2017
// Author:      Michael Toner
// Lab Section: 337-05
// Version:     1.0  Initial Design Entry
// Description: Helper Test Bench Tasks
task send_bit;
begin
end
endtask
