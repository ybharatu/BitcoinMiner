// $Id: $
// File name:   HM_timer.sv
// Created:     11/15/2017
// Author:      Michael Toner
// Lab Section: 337-05
// Version:     1.0  Initial Design Entry
// Description: Flex Counter Wrapper for Hashing Module
