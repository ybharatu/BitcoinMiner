// $Id: $
// File name:   main_controller.sv
// Created:     12/5/2017
// Author:      Yashwanth Bharatula
// Lab Section: 337-05
// Version:     1.0  Initial Design Entry
// Description: Main State Machine
module main_controller
(
	input host_ready,
	input rcv_error,
	output quit_hash,
)


endmodule
